`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////
// Engineer: Bryce Melander
// Company: Cal Poly
//
// Create Date: Dec-18-2023
// Module Name: CSR
// Target Devices: OTTER MCU on Basys3
// Description: 
//
// Dependencies:
//
// Revisions:
//  * 0.01 - File Created
//
// Copyright (c) 2023 by Bryce Melander under MIT License. All rights
// reserved, see http://opensource.org/licenses/MIT for more details.
//////////////////////////////////////////////////////////////////////////////

module CSR (

    );

    initial begin

    end

    always_comb begin

    end

endmodule

// End of File //